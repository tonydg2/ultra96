// for verifying 'axis_stim_syn' only. 

`timescale 1ns / 1ps  // <time_unit>/<time_precision>
  // time_unit: measurement of delays / simulation time (#10 = 10<time_unit>)
  // time_precision: how delay values are rounded before being used in simulation (degree of accuracy of the time unit)

//-------------------------------------------------------------------------------------------------
//
//-------------------------------------------------------------------------------------------------

module led_cnt_tb ;

  logic clk=0, rstn=0, rst;

  //always #2 clk = ~clk; // 250mhz period = 4ns, invert every 2ns
  always #5 clk = ~clk; // 100mhz 

  initial begin
    rstn <= 0;
    #20;
    rstn <= 1;
  end
  assign rst = !rstn;


//-------------------------------------------------------------------------------------------------
//
//-------------------------------------------------------------------------------------------------
//  led_cnt led_cnt(
//    .rst        (rst),
//    .clk100     (clk),
//    .div_i      (5'h1),
//    .wren_i     ('0),
//    .int_clr_i  ('0),
//    .int_cnt_o  (),
//    .led_o      (),
//    .led_int_o  ()
//  );

led_cnt_vhd08 led_cnt_vhd08_inst(
  .rst        (rst),
  .clk        (clk),
  .div_i      (5'h1),
  .wren_i     ('0),
  .led_o      ()
);



endmodule